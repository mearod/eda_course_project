Testbench 1 for homework 4
* For EDA Course 2024

Vin n1 0 10
R1 n1 n2 1
R2 n2 0 4

.dc Vin 10 10 1
.print dc v(n2)

.options NODE

.end
