netlist example

* this is a line of comment

RZjL0 aasd0 0 40
R3 1 2 6k
R4 2 0 0.1

*.op
*.print op v(2)

* Is 0 2 10

.end
